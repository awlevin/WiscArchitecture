module EX_Register();//(clk,rst_n,ALUSrc_in,ALUOp_in,ALUSrc_out,ALUOp_out);
//input clk,rst_n
endmodule

module M_Register();

endmodule

module WB_Register();

endmodule
