module PipelineStages(clk,rst_n);

endmodule

module Fetch();

endmodule

module Decode();

endmodule

module Execute();

endmodule

module Memory();

endmodule

module WriteBack();

endmodule



